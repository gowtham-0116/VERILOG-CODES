module tb;
  reg sel0,sel1;
  reg i0,i1,i2,i3;
  wire y;
   
  mux_3_1 mux(sel0,sel1,i0,i1,i2,i3,y);
  
  initial begin
    $monitor("At time %0t : sel0=%0b,sel1=%0b,i0=%0b,i1=%0b,i2=%0b,i3=%0b,y=%0b",$time , sel0,sel1,i0,i1,i2,i3,y);
    {i3,i2,i1,i0} = 4'h5;

    repeat(8) begin
      {sel0, sel1} = $random;
      #5;
      
      
    end
  end 
endmodule
